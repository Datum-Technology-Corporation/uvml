// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_ST_CHKR_SV__
`define __UVME_ST_CHKR_SV__


/**
 * TODO Describe uvme_st_chkr
 */
module uvme_st_chkr (
      uvma_if  tx_if,
      uvma_if  rx_if
);
   
   // TODO Add assertions to uvme_st_chkr
   
endmodule : uvme_st_chkr


`endif // __UVME_ST_CHKR_SV__
