// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_ST_DUT_CHKR_SV__
`define __UVMT_ST_DUT_CHKR_SV__


/**
 * Module encapsulating assertions for Moore.io UVM Extension LIbrary VIP
 * Self-Testing DUT wrapper (uvmt_st_dut_wrap).
 */
module uvmt_st_dut_chkr(
   uvma_if  tx_if,
   uvma_if  rx_if
);
   
   `pragma protect begin
   
   // TODO Add assertions to uvmt_st_dut_chkr
   
   `pragma protect end
   
endmodule : uvmt_st_dut_chkr


`endif // __UVMT_ST_DUT_CHKR_SV__
