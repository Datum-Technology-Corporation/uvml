// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_ST_IF_CHKR_SV__
`define __UVMA_ST_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_st_if.
 */
module uvma_st_if_chkr(
   uvma_st_if  st_if
);
   
   // TODO Add assertions to uvma_st_if_chkr
   
endmodule : uvma_st_if_chkr


`endif // __UVMA_ST_IF_CHKR_SV__
